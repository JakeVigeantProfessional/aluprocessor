module bit_inverter(data,invertedData);
    input [31:0] data;
    output [31:0] invertedData;
    not not0(invertedData[0], data[0]);
    not not1(invertedData[1], data[1]);
    not not2(invertedData[2], data[2]);
not not3(invertedData[3], data[3]);
not not4(invertedData[4], data[4]);
not not5(invertedData[5], data[5]);
not not6(invertedData[6], data[6]);
not not7(invertedData[7], data[7]);
not not8(invertedData[8], data[8]);
not not9(invertedData[9], data[9]);
not not10(invertedData[10], data[10]);
not not11(invertedData[11], data[11]);
not not12(invertedData[12], data[12]);
not not13(invertedData[13], data[13]);
not not14(invertedData[14], data[14]);
not not15(invertedData[15], data[15]);
not not16(invertedData[16], data[16]);
not not17(invertedData[17], data[17]);
not not18(invertedData[18], data[18]);
not not19(invertedData[19], data[19]);
not not20(invertedData[20], data[20]);
not not21(invertedData[21], data[21]);
not not22(invertedData[22], data[22]);
not not23(invertedData[23], data[23]);
not not24(invertedData[24], data[24]);
not not25(invertedData[25], data[25]);
not not26(invertedData[26], data[26]);
not not27(invertedData[27], data[27]);
not not28(invertedData[28], data[28]);
not not29(invertedData[29], data[29]);
not not30(invertedData[30], data[30]);
not not31(invertedData[31], data[31]);
endmodule